module top;
    integer z;
    initial
        for (integer i; i < 10; i = i + 1)
            z = i;
endmodule
