module testcase;
    wire [3:0] #1 a = 4'b0000;
endmodule
