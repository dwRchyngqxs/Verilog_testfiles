module top;
    reg [2:0] x;
    reg [2:0] x [0:0];
endmodule
