module opt_expr_sub_test4(input [3:0] i, output [8:0] o);
    assign o = 5'b00010 - i;
endmodule
