module top;
    reg [2:0] x [0:0];
    reg [2:0] x;
endmodule
