module top;
    initial begin
        integer x;
    end
endmodule
