module top;
    integer z;
    initial
        for (integer i = 1; i < 10; i = i + 1)
            z = i;
endmodule
