module top;
initial
    begin
        $display("HI");
    end : incorrect_name
endmodule
