module top; wire [7:0] a = (-1)'(a); endmodule
