module foo;

	genvar a;
	for (a = 0; a < 10; a++) begin : a
	end : a
endmodule
