module Example #(
    parameter X, Y
);
endmodule
module top;
    Example #(1) e();
endmodule
