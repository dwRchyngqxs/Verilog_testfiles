module Example #(
    parameter X, Y
);
endmodule
module top;
    Example e();
endmodule
