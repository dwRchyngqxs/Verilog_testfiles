module Task_Test_Top
(
);

    task SomeTaskName(a)
    endtask

endmodule
