module sub (input i, output o);
parameter _TECHMAP_CELLNAME_ = "";
namedsub #(.name(_TECHMAP_CELLNAME_)) _TECHMAP_REPLACE_ (i, o);
endmodule
