module Module #(
    parameter X
);
endmodule
