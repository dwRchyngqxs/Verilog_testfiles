module top (clk, reset, cnt);

input		clk;
input		reset;
output	[7:0]	cnt;

reg	[7:0]	cnt;

endmodule
