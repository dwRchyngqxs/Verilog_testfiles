module test_signed();
parameter logic signed [7:0] a = 0;
parameter logic unsigned [7:0] b = 0;

endmodule
