module top(input [-128:-65] a);
endmodule
