module top(input i, output o);
wire j;
sub s0(i, o, j);
endmodule
