module top(input i, output o, p);
assign o = i;
endmodule
