module m (input i, output o);
wire [1023:0] _TECHMAP_DO_00_ = "CONSTMAP; ";
endmodule
