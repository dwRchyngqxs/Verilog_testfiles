module Example #(
    parameter X
);
endmodule
module top;
    Example e();
endmodule
