module top;
    wire x;
    assign x = 1;
    localparam x = 2;
endmodule
