package correct_name;
localparam X = 1;
endpackage : incorrect_name
