module Module;
    localparam X = 1;
endmodule
