module top2;
	localparam a = 12'h4 /*foo*/'b0;
endmodule
