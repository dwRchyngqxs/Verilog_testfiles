module top(input i, output o);
assign o = i;
endmodule
