module test_signed();
parameter integer signed  a = 0;
parameter integer unsigned  b = 0;

endmodule
