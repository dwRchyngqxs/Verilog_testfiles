module mod;
endmodule
module top;
    reg [2:0] x [0:0];
    mod x();
endmodule
