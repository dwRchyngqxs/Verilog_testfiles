module sub(input i, output o, input j);
wire _TECHMAP_REPLACE_.asdf = i ;
barfoo _TECHMAP_REPLACE_.blah (i, o, j);
endmodule
