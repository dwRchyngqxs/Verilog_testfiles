module top(output o);
m m (.o(o), .i(o));
endmodule
