typedef logic T;
typedef T [3:0] S;
