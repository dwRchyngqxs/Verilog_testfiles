module top;
    initial begin : blk
        integer x;
    end
endmodule
