module sub(input i, output o, (* techmap_autopurge *) input j);
foobar f(i, o, j);
endmodule
