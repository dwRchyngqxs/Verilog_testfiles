module gate(input clk, output [32:0] o, p, q, r, s, t, u);
assign o = 'bx;
assign p = 1'bx;
assign q = 'bz;
assign r = 1'bz;
assign s = 1'b0;
assign t = 'b1;
assign u = -'sb1;
endmodule
