(* src = "\042 \057 \134 \010 \014 \012 \015 \011 \025 \033" *)
module foo;
endmodule
