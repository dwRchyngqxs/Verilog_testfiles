module test_logic_param();
parameter logic                 a = 0;
parameter logic [31:0]          e = 0;
parameter logic signed          b = 0;
parameter logic unsigned        c = 0;
parameter logic unsigned [31:0] d = 0;
endmodule
