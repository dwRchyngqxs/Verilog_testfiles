module test_integer_real();
parameter integer real a = 0;
endmodule
