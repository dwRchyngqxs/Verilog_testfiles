module top; wire [7:0] a = 0'(a); endmodule
