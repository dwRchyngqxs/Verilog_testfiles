module top;
    function automatic integer f;
        input [1:0] inp;
        integer inp;
        f = inp;
    endfunction
    integer x;
    initial x = f(0);
endmodule
