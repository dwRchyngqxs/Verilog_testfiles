module top(input i, output o);
sub s0(i, o);
endmodule
