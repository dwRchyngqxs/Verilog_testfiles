// megafunction wizard: %ALTMULT_ACCUM (MAC)%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altmult_add 

// ============================================================
// File Name: scanout_chain_megafn.v
// Megafunction Name(s):
// 			altmult_add
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Build 178 05/31/2012 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2012 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module scanout_chain_megafn (
	clock0,
	dataa_0,
	datab_0,
	datab_1,
	datab_2,
	datab_3,
	result,
	shiftouta);

	input	  clock0;
	input	[17:0]  dataa_0;
	input	[17:0]  datab_0;
	input	[17:0]  datab_1;
	input	[17:0]  datab_2;
	input	[17:0]  datab_3;
	output	[43:0]  result;
	output	[17:0]  shiftouta;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  clock0;
	tri0	[17:0]  dataa_0;
	tri0	[17:0]  datab_0;
	tri0	[17:0]  datab_1;
	tri0	[17:0]  datab_2;
	tri0	[17:0]  datab_3;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACCUM_DIRECTION STRING "Add"
// Retrieval info: PRIVATE: ACCUM_SLOAD NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPELINE_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPELINE_REG NUMERIC "1"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPELINE_REG_INDEX NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ACCUM_SLOAD_REG NUMERIC "1"
// Retrieval info: PRIVATE: ACCUM_SLOAD_REG_INDEX NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_PIPELINE_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_PIPELINE_REG NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_REG NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB1_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB1_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB1_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB1_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB1_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ADDNSUB1_REG STRING "1"
// Retrieval info: PRIVATE: ADDNSUB3_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB3_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB3_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB3_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB3_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ADDNSUB3_REG STRING "1"
// Retrieval info: PRIVATE: ADD_ENABLE NUMERIC "0"
// Retrieval info: PRIVATE: ALL_REG_ACLR NUMERIC "0"
// Retrieval info: PRIVATE: A_ACLR_SRC_MULT0 NUMERIC "3"
// Retrieval info: PRIVATE: A_CLK_SRC_MULT0 NUMERIC "0"
// Retrieval info: PRIVATE: B_ACLR_SRC_MULT0 NUMERIC "3"
// Retrieval info: PRIVATE: B_CLK_SRC_MULT0 NUMERIC "0"
// Retrieval info: PRIVATE: CHAINOUT_OUTPUT_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: CHAINOUT_OUTPUT_REG STRING "0"
// Retrieval info: PRIVATE: CHAINOUT_OUTPUT_REGISTER NUMERIC "0"
// Retrieval info: PRIVATE: CHAINOUT_OUTPUT_REGISTERED NUMERIC "0"
// Retrieval info: PRIVATE: CHAS_ZERO_CHAINOUT NUMERIC "0"
// Retrieval info: PRIVATE: EXTRA_MULTIPLIER_LATENCY NUMERIC "0"
// Retrieval info: PRIVATE: HAS_ACCUMULATOR NUMERIC "1"
// Retrieval info: PRIVATE: HAS_ACUMM_SLOAD NUMERIC "0"
// Retrieval info: PRIVATE: HAS_CHAININ_PORT NUMERIC "0"
// Retrieval info: PRIVATE: HAS_CHAINOUT_ADDER NUMERIC "0"
// Retrieval info: PRIVATE: HAS_LOOPBACK NUMERIC "0"
// Retrieval info: PRIVATE: HAS_MAC STRING "1"
// Retrieval info: PRIVATE: HAS_SAT_ROUND STRING "1"
// Retrieval info: PRIVATE: HAS_ZERO_LOOPBACK NUMERIC "0"
// Retrieval info: PRIVATE: IMPL_STYLE_DEDICATED NUMERIC "1"
// Retrieval info: PRIVATE: IMPL_STYLE_DEFAULT NUMERIC "0"
// Retrieval info: PRIVATE: IMPL_STYLE_LCELL NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: PRIVATE: MULT_LATENCY NUMERIC "0"
// Retrieval info: PRIVATE: MULT_REGA0 NUMERIC "1"
// Retrieval info: PRIVATE: MULT_REGB0 NUMERIC "1"
// Retrieval info: PRIVATE: MULT_REGOUT0 NUMERIC "1"
// Retrieval info: PRIVATE: NUM_MULT STRING "4"
// Retrieval info: PRIVATE: OP1 STRING "Add"
// Retrieval info: PRIVATE: OP3 STRING "Add"
// Retrieval info: PRIVATE: OUTPUT_EXTRA_LAT NUMERIC "0"
// Retrieval info: PRIVATE: OUTPUT_REG_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: OUTPUT_REG_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: OVERFLOW NUMERIC "0"
// Retrieval info: PRIVATE: Q_ACLR_SRC_MULT0 NUMERIC "3"
// Retrieval info: PRIVATE: Q_CLK_SRC_MULT0 NUMERIC "0"
// Retrieval info: PRIVATE: REG_OUT NUMERIC "1"
// Retrieval info: PRIVATE: RNFORMAT STRING "44"
// Retrieval info: PRIVATE: ROTATE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROTATE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROTATE_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROTATE_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROTATE_OUT_REG STRING "1"
// Retrieval info: PRIVATE: ROTATE_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROTATE_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROTATE_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ROTATE_REG STRING "1"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_MODE STRING "Disabled"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_OUT_REG STRING "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_REG STRING "1"
// Retrieval info: PRIVATE: ROUND3_FRAC_WIDTH NUMERIC "23"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_CHAINOUT_TYPE STRING "Nearest Integer"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_MODE STRING "Disabled"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_REG STRING "1"
// Retrieval info: PRIVATE: RQFORMAT STRING "Q1.30"
// Retrieval info: PRIVATE: RTS_WIDTH STRING "44"
// Retrieval info: PRIVATE: SAME_CONFIG NUMERIC "1"
// Retrieval info: PRIVATE: SAME_CONTROL_SRC_A0 NUMERIC "1"
// Retrieval info: PRIVATE: SAME_CONTROL_SRC_B0 NUMERIC "1"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_MODE STRING "Enabled"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_REG STRING "1"
// Retrieval info: PRIVATE: SAT3_FRAC_WIDTH NUMERIC "1"
// Retrieval info: PRIVATE: SAT3_OUTPUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_OUTPUT_CHAINOUT_TYPE STRING "Symmetric"
// Retrieval info: PRIVATE: SAT3_OUTPUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_OUTPUT_MODE STRING "Enabled"
// Retrieval info: PRIVATE: SAT3_OUTPUT_OVERFLOW NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_OUTPUT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_OUTPUT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_OUTPUT_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: SAT3_OUTPUT_REG STRING "1"
// Retrieval info: PRIVATE: SCANOUTA NUMERIC "1"
// Retrieval info: PRIVATE: SCANOUTB NUMERIC "0"
// Retrieval info: PRIVATE: SHIFTOUTA_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFTOUTA_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFTOUTA_REG STRING "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFT_RIGHT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFT_RIGHT_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_OUT_REG STRING "1"
// Retrieval info: PRIVATE: SHIFT_RIGHT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFT_RIGHT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: SHIFT_RIGHT_REG STRING "1"
// Retrieval info: PRIVATE: SHIFT_ROTATE_MODE STRING "None"
// Retrieval info: PRIVATE: SIGNA STRING "SIGNED"
// Retrieval info: PRIVATE: SIGNA_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNA_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNA_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNA_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNA_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: SIGNA_REG STRING "1"
// Retrieval info: PRIVATE: SIGNB STRING "SIGNED"
// Retrieval info: PRIVATE: SIGNB_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNB_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNB_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNB_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNB_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: SIGNB_REG STRING "1"
// Retrieval info: PRIVATE: SRCA0 STRING "Shiftin input"
// Retrieval info: PRIVATE: SRCB0 STRING "Multiplier input"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: WIDTHA STRING "18"
// Retrieval info: PRIVATE: WIDTHB STRING "18"
// Retrieval info: PRIVATE: WIDTH_UPPER_DATA NUMERIC "1"
// Retrieval info: PRIVATE: ZERO_CHAINOUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ZERO_CHAINOUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_CHAINOUT_REG STRING "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_OUT_REG STRING "1"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_REG STRING "1"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: ACCUMULATOR STRING "YES"
// Retrieval info: CONSTANT: ACCUM_DIRECTION STRING "ADD"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_ACLR1 STRING "UNUSED"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_ACLR3 STRING "UNUSED"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_ACLR1 STRING "UNUSED"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_ACLR3 STRING "UNUSED"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_REGISTER1 STRING "CLOCK0"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_REGISTER3 STRING "CLOCK0"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_REGISTER1 STRING "CLOCK0"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_REGISTER3 STRING "CLOCK0"
// Retrieval info: CONSTANT: CHAINOUT_ADDER STRING "NO"
// Retrieval info: CONSTANT: CHAINOUT_REGISTER STRING "UNREGISTERED"
// Retrieval info: CONSTANT: DEDICATED_MULTIPLIER_CIRCUITRY STRING "YES"
// Retrieval info: CONSTANT: INPUT_ACLR_A0 STRING "UNUSED"
// Retrieval info: CONSTANT: INPUT_ACLR_A1 STRING "UNUSED"
// Retrieval info: CONSTANT: INPUT_ACLR_A2 STRING "UNUSED"
// Retrieval info: CONSTANT: INPUT_ACLR_A3 STRING "UNUSED"
// Retrieval info: CONSTANT: INPUT_ACLR_B0 STRING "UNUSED"
// Retrieval info: CONSTANT: INPUT_ACLR_B1 STRING "UNUSED"
// Retrieval info: CONSTANT: INPUT_ACLR_B2 STRING "UNUSED"
// Retrieval info: CONSTANT: INPUT_ACLR_B3 STRING "UNUSED"
// Retrieval info: CONSTANT: INPUT_REGISTER_A0 STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_REGISTER_A1 STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_REGISTER_A2 STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_REGISTER_A3 STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_REGISTER_B0 STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_REGISTER_B1 STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_REGISTER_B2 STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_REGISTER_B3 STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_SOURCE_A0 STRING "DATAA"
// Retrieval info: CONSTANT: INPUT_SOURCE_A1 STRING "SCANA"
// Retrieval info: CONSTANT: INPUT_SOURCE_A2 STRING "SCANA"
// Retrieval info: CONSTANT: INPUT_SOURCE_A3 STRING "SCANA"
// Retrieval info: CONSTANT: INPUT_SOURCE_B0 STRING "DATAB"
// Retrieval info: CONSTANT: INPUT_SOURCE_B1 STRING "DATAB"
// Retrieval info: CONSTANT: INPUT_SOURCE_B2 STRING "DATAB"
// Retrieval info: CONSTANT: INPUT_SOURCE_B3 STRING "DATAB"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altmult_add"
// Retrieval info: CONSTANT: MULTIPLIER1_DIRECTION STRING "ADD"
// Retrieval info: CONSTANT: MULTIPLIER3_DIRECTION STRING "ADD"
// Retrieval info: CONSTANT: MULTIPLIER_ACLR0 STRING "UNUSED"
// Retrieval info: CONSTANT: MULTIPLIER_ACLR1 STRING "UNUSED"
// Retrieval info: CONSTANT: MULTIPLIER_ACLR2 STRING "UNUSED"
// Retrieval info: CONSTANT: MULTIPLIER_ACLR3 STRING "UNUSED"
// Retrieval info: CONSTANT: MULTIPLIER_REGISTER0 STRING "CLOCK0"
// Retrieval info: CONSTANT: MULTIPLIER_REGISTER1 STRING "CLOCK0"
// Retrieval info: CONSTANT: MULTIPLIER_REGISTER2 STRING "CLOCK0"
// Retrieval info: CONSTANT: MULTIPLIER_REGISTER3 STRING "CLOCK0"
// Retrieval info: CONSTANT: NUMBER_OF_MULTIPLIERS NUMERIC "4"
// Retrieval info: CONSTANT: OUTPUT_ACLR STRING "UNUSED"
// Retrieval info: CONSTANT: OUTPUT_REGISTER STRING "CLOCK0"
// Retrieval info: CONSTANT: OUTPUT_ROUND_TYPE STRING "NEAREST_INTEGER"
// Retrieval info: CONSTANT: OUTPUT_SATURATE_ACLR STRING "UNUSED"
// Retrieval info: CONSTANT: OUTPUT_SATURATE_PIPELINE_ACLR STRING "UNUSED"
// Retrieval info: CONSTANT: OUTPUT_SATURATE_PIPELINE_REGISTER STRING "CLOCK0"
// Retrieval info: CONSTANT: OUTPUT_SATURATE_REGISTER STRING "CLOCK0"
// Retrieval info: CONSTANT: OUTPUT_SATURATE_TYPE STRING "SYMMETRIC"
// Retrieval info: CONSTANT: OUTPUT_SATURATION STRING "YES"
// Retrieval info: CONSTANT: PORT_ADDNSUB1 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_ADDNSUB3 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SIGNA STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SIGNB STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: REPRESENTATION_A STRING "SIGNED"
// Retrieval info: CONSTANT: REPRESENTATION_B STRING "SIGNED"
// Retrieval info: CONSTANT: SCANOUTA_REGISTER STRING "UNREGISTERED"
// Retrieval info: CONSTANT: SIGNED_ACLR_A STRING "UNUSED"
// Retrieval info: CONSTANT: SIGNED_ACLR_B STRING "UNUSED"
// Retrieval info: CONSTANT: SIGNED_PIPELINE_ACLR_A STRING "UNUSED"
// Retrieval info: CONSTANT: SIGNED_PIPELINE_ACLR_B STRING "UNUSED"
// Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_A STRING "CLOCK0"
// Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_B STRING "CLOCK0"
// Retrieval info: CONSTANT: SIGNED_REGISTER_A STRING "CLOCK0"
// Retrieval info: CONSTANT: SIGNED_REGISTER_B STRING "CLOCK0"
// Retrieval info: CONSTANT: WIDTH_A NUMERIC "18"
// Retrieval info: CONSTANT: WIDTH_B NUMERIC "18"
// Retrieval info: CONSTANT: WIDTH_CHAININ NUMERIC "1"
// Retrieval info: CONSTANT: WIDTH_MSB NUMERIC "44"
// Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "44"
// Retrieval info: CONSTANT: WIDTH_SATURATE_SIGN NUMERIC "1"
// Retrieval info: CONSTANT: ZERO_CHAINOUT_OUTPUT_ACLR STRING "UNUSED"
// Retrieval info: CONSTANT: ZERO_CHAINOUT_OUTPUT_REGISTER STRING "CLOCK0"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_ACLR STRING "UNUSED"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_OUTPUT_ACLR STRING "UNUSED"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_OUTPUT_REGISTER STRING "CLOCK0"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_PIPELINE_ACLR STRING "UNUSED"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_PIPELINE_REGISTER STRING "CLOCK0"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_REGISTER STRING "CLOCK0"
// Retrieval info: USED_PORT: clock0 0 0 0 0 INPUT VCC "clock0"
// Retrieval info: USED_PORT: dataa_0 0 0 18 0 INPUT GND "dataa_0[17..0]"
// Retrieval info: USED_PORT: datab_0 0 0 18 0 INPUT GND "datab_0[17..0]"
// Retrieval info: USED_PORT: datab_1 0 0 18 0 INPUT GND "datab_1[17..0]"
// Retrieval info: USED_PORT: datab_2 0 0 18 0 INPUT GND "datab_2[17..0]"
// Retrieval info: USED_PORT: datab_3 0 0 18 0 INPUT GND "datab_3[17..0]"
// Retrieval info: USED_PORT: result 0 0 44 0 OUTPUT GND "result[43..0]"
// Retrieval info: USED_PORT: shiftouta 0 0 18 0 OUTPUT GND "shiftouta[17..0]"
// Retrieval info: CONNECT: @clock0 0 0 0 0 clock0 0 0 0 0
// Retrieval info: CONNECT: @dataa 0 0 18 18 GND 0 0 18 0
// Retrieval info: CONNECT: @dataa 0 0 18 36 GND 0 0 18 0
// Retrieval info: CONNECT: @dataa 0 0 18 54 GND 0 0 18 0
// Retrieval info: CONNECT: @dataa 0 0 18 0 dataa_0 0 0 18 0
// Retrieval info: CONNECT: @datab 0 0 18 0 datab_0 0 0 18 0
// Retrieval info: CONNECT: @datab 0 0 18 18 datab_1 0 0 18 0
// Retrieval info: CONNECT: @datab 0 0 18 36 datab_2 0 0 18 0
// Retrieval info: CONNECT: @datab 0 0 18 54 datab_3 0 0 18 0
// Retrieval info: CONNECT: result 0 0 44 0 @result 0 0 44 0
// Retrieval info: CONNECT: shiftouta 0 0 18 0 @scanouta 0 0 18 0
// Retrieval info: GEN_FILE: TYPE_NORMAL scanout_chain_megafn.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL scanout_chain_megafn.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL scanout_chain_megafn.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL scanout_chain_megafn.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL scanout_chain_megafn_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL scanout_chain_megafn_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
