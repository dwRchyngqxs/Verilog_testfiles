module top;
initial
    begin : correct_name
        $display("HI");
    end : incorrect_name
endmodule
