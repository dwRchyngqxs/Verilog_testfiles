module top; wire [7:0] a, b = (a)'(0); endmodule
