module top;
if (1)
    begin : correct_name
        initial $display("HI");
    end : incorrect_name
endmodule
