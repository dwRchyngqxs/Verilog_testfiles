module DFF(input D, C, output Q);
endmodule
