module top;
    for (genvar i = 1; i < 10; i = i + 1)
        wire x;
endmodule
