module test_signed();
parameter signed integer a = 0;
parameter unsigned integer b = 0;

endmodule
