module sub(input i, output o, (* techmap_autopurge *) input [1:0] j);
foobar f(i, o, j);
endmodule
