module Example #(
    parameter X, Y
);
endmodule
module top;
    Example #(.Y(1)) e();
endmodule
