module correct_name;
localparam X = 1;
endmodule : incorrect_name
