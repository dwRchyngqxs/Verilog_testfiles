module correct_name;
localparam X = 1;
endmodule : correct_name
