module gold(input i, output o);
assign o = 1'bx ~^ i;
endmodule
