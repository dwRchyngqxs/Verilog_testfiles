module foo3;

	genvar a;
	for (a = 0; a < 10; a++) begin : a
	end : b
endmodule
