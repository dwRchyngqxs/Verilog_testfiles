module test;
    reg q;
    initial #(1) q = 1;
endmodule
