module top;
    for (genvar i; i < 10; i = i + 1)
        wire x;
endmodule
