package correct_name;
localparam X = 1;
endpackage : correct_name
