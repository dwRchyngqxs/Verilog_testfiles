module top();
    wire a, b, c;
endmodule
