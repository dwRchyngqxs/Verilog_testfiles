parameter Q = 1;
