module test_integer_range();
parameter integer [31:0] a = 0;
endmodule
