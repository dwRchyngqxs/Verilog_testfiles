module Module #(
    localparam X
);
endmodule
