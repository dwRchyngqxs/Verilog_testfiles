module top;
if (1)
    begin
        initial $display("HI");
    end : incorrect_name
endmodule
